library verilog;
use verilog.vl_types.all;
entity Sequence_Detector_vlg_vec_tst is
end Sequence_Detector_vlg_vec_tst;
