library verilog;
use verilog.vl_types.all;
entity TIMER_vlg_vec_tst is
end TIMER_vlg_vec_tst;
