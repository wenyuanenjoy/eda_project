library verilog;
use verilog.vl_types.all;
entity APB_Slave_vlg_vec_tst is
end APB_Slave_vlg_vec_tst;
